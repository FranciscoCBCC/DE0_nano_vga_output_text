LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
 
ENTITY PixelGen IS
	PORT(
		RESET : IN STD_LOGIC; -- Entrada para reiniciar o estado do controlador
		F_CLOCK : IN STD_LOGIC; -- Entrada de clock (50 MHz)
		F_ON : IN STD_LOGIC; --Indica a região ativa do frame
		F_ROW : IN STD_LOGIC_VECTOR(9 DOWNTO 0); -- Índice da linha que está sendo processada
		F_COLUMN : IN STD_LOGIC_VECTOR(10 DOWNTO 0); -- Índice da coluna que está sendo processada
		R_OUT : OUT STD_LOGIC; -- Componente R
		G_OUT : OUT STD_LOGIC; -- Componente G
		B_OUT : OUT STD_LOGIC -- Componente B
	);
 
END ENTITY PixelGen;
 
ARCHITECTURE arch OF PixelGen IS
 
 COMPONENT font_rom IS
	port(
		clk: in std_logic;
		addr: in std_logic_vector(10 downto 0);
		data: out std_logic_vector(7 downto 0)
	);
 END COMPONENT font_rom;
 
 --Coordenadas X e Y do pixel atual
   SIGNAL pix_x, pix_y: UNSIGNED(9 DOWNTO 0);
 
 --Endereço que será acessado na memória de caracteres
   SIGNAL rom_addr: STD_LOGIC_VECTOR(10 DOWNTO 0);
 
 --Código ASCII do caractere atual (parte do endereço)
   SIGNAL char_addr: STD_LOGIC_VECTOR(6 DOWNTO 0);
 
 --Parte do caractere (0~15) que está sendo exibida na linha atual Y
   SIGNAL row_addr: STD_LOGIC_VECTOR(3 DOWNTO 0);
 
 --Pixel relativo a coordenada X atual
   SIGNAL bit_addr: STD_LOGIC_VECTOR(2 DOWNTO 0);
 
 --Conteúdo armazenado no endereço indicado por 'rom_addr'
   SIGNAL font_word: STD_LOGIC_VECTOR(7 DOWNTO 0);
 
 --Valor do bit 'bit_addr' na palavra 'font_word'
   SIGNAL font_bit: STD_LOGIC;
 
 --Valor das componentes rgb
   SIGNAL font_rgb: STD_LOGIC_VECTOR(2 DOWNTO 0);
 
 --Flag que indica se a frase deve ser exibida
   SIGNAL txt_on: STD_LOGIC;
 
BEGIN
 
 -- Coordenadas XY atuais
 pix_x <= UNSIGNED(F_COLUMN(9 DOWNTO 0));
 pix_y <= UNSIGNED(F_ROW);
 
 -- Memória dos caracteres
 font_unit: font_rom PORT MAP(clk=>not F_CLOCK, addr=>rom_addr, data=>font_word);
 
 -- Determinação do endereço que será acessado
 row_addr <= STD_LOGIC_VECTOR(pix_y(3 DOWNTO 0));
 rom_addr <= char_addr & row_addr;
 
   txt_on <= '1' WHEN (pix_x >= 320 AND pix_x <= 455) AND (pix_y >= 292 AND pix_y <= 305) ELSE
              '0';
   
   WITH pix_x(7 DOWNTO 3) SELECT
     char_addr <=
 "1100110" WHEN "01000", -- f
 "1110010" WHEN "01001", -- r
 "1100001" WHEN "01010", -- a
 "1101110" WHEN "01011", -- n
 "1100011" WHEN "01100", -- c
 "1101001" WHEN "01101", -- i
 "1110011" WHEN "01110", -- s
 "1100011" WHEN "01111", -- c
 "1101111" WHEN "10000", -- o
 "0000000" WHEN "10001", --
 "0000000" WHEN OTHERS;
   
 
 bit_addr <= NOT STD_LOGIC_VECTOR(pix_x(2 DOWNTO 0));
 font_bit <= font_word(to_integer(UNSIGNED( bit_addr))); 
 
 font_rgb <="111" WHEN font_bit='1' ELSE "000";
 
 PROCESS(F_ON,font_rgb,txt_on)
 BEGIN
 
 IF F_ON ='0' or txt_on='0' THEN
 R_OUT <= '0';
 G_OUT <= '0';
 B_OUT <= '0';
 ELSE
 R_OUT <= font_rgb(0);
 G_OUT <= font_rgb(1);
 B_OUT <= font_rgb(2); 
 END IF;
 END PROCESS; 
 
END ARCHITECTURE arch;